LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY leddec IS
	PORT (
		dig : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		data : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		displays : OUT STD_LOGIC_VECTOR (41 DOWNTO 0)
		--seg : OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
	);
END leddec;

ARCHITECTURE Behavioral OF leddec IS
	SIGNAL seg : STD_LOGIC_VECTOR (6 DOWNTO 0);
BEGIN

	-- Turn on segments corresponding to 4-bit data word
	seg <= "0000001" WHEN data = "0000" ELSE --0
	       "1001111" WHEN data = "0001" ELSE --1
	       "0010010" WHEN data = "0010" ELSE --2
	       "0000110" WHEN data = "0011" ELSE --3
	       "1001100" WHEN data = "0100" ELSE --4
	       "0100100" WHEN data = "0101" ELSE --5
	       "0100000" WHEN data = "0110" ELSE --6
	       "0001111" WHEN data = "0111" ELSE --7
	       "0000000" WHEN data = "1000" ELSE --8
	       "0000100" WHEN data = "1001" ELSE --9
	       "0001000" WHEN data = "1010" ELSE --A
	       "1100000" WHEN data = "1011" ELSE --B
	       "0110001" WHEN data = "1100" ELSE --C
	       "1000010" WHEN data = "1101" ELSE --D
	       "0110000" WHEN data = "1110" ELSE --E
	       "0111000" WHEN data = "1111" ELSE --F
	       "1111111";
	-- Turn on anode of 7-segment display addressed by 2-bit digit selector dig for Nexys board
	--anode <= "1110" WHEN dig = "00" ELSE --0
	--         "1101" WHEN dig = "01" ELSE --1
	--         "1011" WHEN dig = "10" ELSE --2
	--         "0111" WHEN dig = "11" ELSE --3
	--         "1111";
	-- Turn on 1 of 6 7-segment display addressed by 3-bit digit selector dig for Terasic DE0-CV
process(dig)
begin
		if (dig = "000") then 
		   displays (41 DOWNTO 35) <= seg;
		elsif (dig = "001") then
			displays (34 DOWNTO 28) <= seg;
		elsif (dig = "010") then
			displays (27 DOWNTO 21) <= seg;
		elsif (dig = "110") then--011 is translated to 110 why? 110 is 011 and 011 is 110?
			displays (20 DOWNTO 14) <= seg;
		elsif (dig = "100") then
			displays (13 DOWNTO 7) <= seg;
		elsif (dig = "101") then
			displays (6 DOWNTO 0) <= seg;
		else 
		end if;
end process;
END Behavioral;
