LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY hexcount IS
	PORT (
		clk_50MHz : IN STD_LOGIC;
		--anode : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		displays : OUT STD_LOGIC_VECTOR (41 DOWNTO 0);
		--seg : OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
		swt: IN STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
END hexcount;

ARCHITECTURE Behavioral OF hexcount IS
	COMPONENT counter IS
		PORT (
			clk : IN STD_LOGIC;
			count : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT leddec IS
		PORT (
			dig : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			data : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			--anode : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			--seg : OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
			displays : OUT STD_LOGIC_VECTOR (41 DOWNTO 0)
		);
	END COMPONENT;
	SIGNAL S : STD_LOGIC_VECTOR (3 DOWNTO 0);
BEGIN
	C1 : counter
	PORT MAP(clk => clk_50MHz, count => S);
	L1 : leddec
	--PORT MAP(dig => "00", data => S, anode => anode, seg => seg);
	PORT MAP(dig => swt, data => S, displays => displays);
END Behavioral;
